module instruction (input [31:0] address,
                       output [31:0] instruction);
    
    reg [31:0] memory [63:0];

    // ADDi $1, R[0], R[6]
    // "000000000001_00000_000_00110_0010000"
    assign memory[0] = 32'b00000000000100000000001100010000;

    // ADDi $0, R[0], R[7]
    // "000000000000_00000_000_00111_0010000"
    assign memory[4] = 32'b00000000000000000000001110010000;

    // ADDi $0, R[6],  R[8]
    // "000000000000_00110_000_01000_0010000"
    assign memory[8] = 32'b00000000000000110000010000010000;

    // ADD R[7], R[6], R[6]
    // "0000000_00111_00110_000_00110_0110000"
    assign memory[12] = 32'b00000000011100110000001100110000;

    // ADDi $0, R[8], R[7]
    // "000000000000_01000_000_00111_0010000"
    assign memory[16] = 32'b00000000000001000000001110010000;

    // JUMP 
    // 111111111111_11111_101_00111_1101100
    assign memory[20] = 32'b11111111111111111101001111101100;

    assign instruction = memory[address];

endmodule

// -- result(1) := "00000000001100110000010000010000";

// -- "000000000000_00000_000_00110_0010000"
// result(0) := "00000000000100000000001100010000";
// -- "000000000001_00000_000_00111_0010000"
// result(1) := "00000000000000000000001110010000";

// -- "000000000000_00110_000_01000_0010000"
// result(2) := "00000000000000110000010000010000";
// -- "0000000_00111_00110_000_00110_0110000"
// result(3) := "00000000011100110000001100110000";
// -- "000000000000_01000_000_00111_0010000"
// result(4) := "00000000000001000000001110010000";

// -- 111111111111_11111_110_00111_1101100
// result(5) := "11111111111111111101001111101100";