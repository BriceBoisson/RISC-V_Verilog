parameter [2:0] LB  = 3'b000;
parameter [2:0] LH  = 3'b001;
parameter [2:0] LW  = 3'b010;
parameter [2:0] LBU = 3'b011;
parameter [2:0] LHU = 3'b100;

parameter [2:0] SB  = 2'b00;
parameter [2:0] SH  = 2'b01;
parameter [2:0] SW  = 2'b10;
