module tb_alu (S);
    output [31:0] S;
endmodule